
package calc_tb_pkg;
  import calculator_pkg::*;
  `include "calc_seq_item.svh"
  `include "calc_driver.svh"
  `include "calc_monitor.svh"
  `include "calc_sequencer.svh"
  `include "calc_sb.svh"

endpackage : calc_tb_pkg


